`define ADDER_WIDTH 32